`default_nettype none
`timescale 1ns/1ns

/* FP32 Divitor Design
*TODO: make a TODO list
*/
module FP32_Div #(
) ()



endmodule